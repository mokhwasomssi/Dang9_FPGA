reg [9:0] deg, Vx, Vy, Dx, Dy, R;

always @(posedge clk or posedge rst)
    if(rst) begin
    end
    else begin
        case(R)
            12 : case(deg)
                0	:	begin	Vx	=	12	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	3	;	Vy	=	12	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	11	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	10	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end
                20	:	begin	Vx	=	4	;	Vy	=	10	;	Dx	=	1	;	Dy	=	-1	;	end
                25	:	begin	Vx	=	11	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	1	;	Vy	=	12	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	11	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	9	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
                45	:	begin	Vx	=	6	;	Vy	=	10	;	Dx	=	1	;	Dy	=	-1	;	end
                50	:	begin	Vx	=	11	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	12	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	12	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	7	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	-1	;	end
                70	:	begin	Vx	=	7	;	Vy	=	9	;	Dx	=	1	;	Dy	=	-1	;	end
                75	:	begin	Vx	=	11	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	2	;	Vy	=	12	;	Dx	=	-1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	12	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	6	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	-1	;	end
                95	:	begin	Vx	=	8	;	Vy	=	8	;	Dx	=	1	;	Dy	=	-1	;	end
                100	:	begin	Vx	=	10	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	3	;	Vy	=	12	;	Dx	=	-1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	12	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	4	;	Vy	=	11	;	Dx	=	-1	;	Dy	=	-1	;	end
                120	:	begin	Vx	=	9	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                125	:	begin	Vx	=	9	;	Vy	=	8	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	5	;	Vy	=	12	;	Dx	=	-1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	12	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                140	:	begin	Vx	=	3	;	Vy	=	11	;	Dx	=	-1	;	Dy	=	-1	;	end
                145	:	begin	Vx	=	10	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                150	:	begin	Vx	=	8	;	Vy	=	9	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	6	;	Vy	=	11	;	Dx	=	-1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	12	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                165	:	begin	Vx	=	1	;	Vy	=	11	;	Dx	=	-1	;	Dy	=	-1	;	end
                170	:	begin	Vx	=	11	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                175	:	begin	Vx	=	7	;	Vy	=	10	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	8	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	12	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	11	;	Dx	=	1	;	Dy	=	-1	;	end
                195	:	begin	Vx	=	11	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                200	:	begin	Vx	=	5	;	Vy	=	11	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	9	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	11	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                215	:	begin	Vx	=	2	;	Vy	=	11	;	Dx	=	1	;	Dy	=	-1	;	end
                220	:	begin	Vx	=	11	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                225	:	begin	Vx	=	4	;	Vy	=	12	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	10	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	10	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                240	:	begin	Vx	=	3	;	Vy	=	11	;	Dx	=	1	;	Dy	=	-1	;	end
                245	:	begin	Vx	=	11	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	2	;	Vy	=	12	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	11	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	9	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
                265	:	begin	Vx	=	5	;	Vy	=	10	;	Dx	=	1	;	Dy	=	-1	;	end
                270	:	begin	Vx	=	11	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	1	;	Vy	=	12	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	12	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	8	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	-1	;	end
                290	:	begin	Vx	=	6	;	Vy	=	9	;	Dx	=	1	;	Dy	=	-1	;	end
                295	:	begin	Vx	=	11	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	1	;	Vy	=	12	;	Dx	=	-1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	12	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	7	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	-1	;	end
                315	:	begin	Vx	=	8	;	Vy	=	8	;	Dx	=	1	;	Dy	=	-1	;	end
                320	:	begin	Vx	=	10	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	2	;	Vy	=	12	;	Dx	=	-1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	12	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	5	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	-1	;	end
                340	:	begin	Vx	=	9	;	Vy	=	7	;	Dx	=	1	;	Dy	=	-1	;	end
                345	:	begin	Vx	=	10	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	4	;	Vy	=	12	;	Dx	=	-1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	12	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	4	;	Vy	=	11	;	Dx	=	-1	;	Dy	=	-1	;	end
            endcase
            11 : case(deg)
                0	:	begin	Vx	=	11	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	3	;	Vy	=	11	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	10	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	9	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end
                20	:	begin	Vx	=	4	;	Vy	=	10	;	Dx	=	1	;	Dy	=	-1	;	end
                25	:	begin	Vx	=	10	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	1	;	Vy	=	11	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	10	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	8	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
                45	:	begin	Vx	=	5	;	Vy	=	9	;	Dx	=	1	;	Dy	=	-1	;	end
                50	:	begin	Vx	=	10	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	11	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	11	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	7	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	-1	;	end
                70	:	begin	Vx	=	6	;	Vy	=	8	;	Dx	=	1	;	Dy	=	-1	;	end
                75	:	begin	Vx	=	10	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	2	;	Vy	=	11	;	Dx	=	-1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	11	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	5	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	-1	;	end
                95	:	begin	Vx	=	8	;	Vy	=	7	;	Dx	=	1	;	Dy	=	-1	;	end
                100	:	begin	Vx	=	9	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	3	;	Vy	=	11	;	Dx	=	-1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	11	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	4	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	-1	;	end
                120	:	begin	Vx	=	8	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                125	:	begin	Vx	=	8	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	5	;	Vy	=	11	;	Dx	=	-1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	11	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                140	:	begin	Vx	=	3	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	-1	;	end
                145	:	begin	Vx	=	9	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                150	:	begin	Vx	=	7	;	Vy	=	8	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	6	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	11	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                165	:	begin	Vx	=	1	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	-1	;	end
                170	:	begin	Vx	=	10	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                175	:	begin	Vx	=	6	;	Vy	=	9	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	7	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	11	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	10	;	Dx	=	1	;	Dy	=	-1	;	end
                195	:	begin	Vx	=	10	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                200	:	begin	Vx	=	5	;	Vy	=	10	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	8	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	10	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                215	:	begin	Vx	=	2	;	Vy	=	10	;	Dx	=	1	;	Dy	=	-1	;	end
                220	:	begin	Vx	=	10	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                225	:	begin	Vx	=	4	;	Vy	=	11	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	9	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	9	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                240	:	begin	Vx	=	3	;	Vy	=	10	;	Dx	=	1	;	Dy	=	-1	;	end
                245	:	begin	Vx	=	10	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	2	;	Vy	=	11	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	10	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	9	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end
                265	:	begin	Vx	=	4	;	Vy	=	9	;	Dx	=	1	;	Dy	=	-1	;	end
                270	:	begin	Vx	=	10	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	1	;	Vy	=	11	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	11	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	7	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
                290	:	begin	Vx	=	6	;	Vy	=	9	;	Dx	=	1	;	Dy	=	-1	;	end
                295	:	begin	Vx	=	10	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	1	;	Vy	=	11	;	Dx	=	-1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	11	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	6	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	-1	;	end
                315	:	begin	Vx	=	7	;	Vy	=	8	;	Dx	=	1	;	Dy	=	-1	;	end
                320	:	begin	Vx	=	9	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	2	;	Vy	=	11	;	Dx	=	-1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	11	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	5	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	-1	;	end
                340	:	begin	Vx	=	8	;	Vy	=	7	;	Dx	=	1	;	Dy	=	-1	;	end
                345	:	begin	Vx	=	9	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	4	;	Vy	=	11	;	Dx	=	-1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	11	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	4	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	-1	;	end

            endcase
            10 : case(deg)
                0	:	begin	Vx	=	10	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	2	;	Vy	=	10	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	9	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	8	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                20	:	begin	Vx	=	4	;	Vy	=	9	;	Dx	=	1	;	Dy	=	-1	;	end
                25	:	begin	Vx	=	9	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	1	;	Vy	=	10	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	10	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	7	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end
                45	:	begin	Vx	=	5	;	Vy	=	8	;	Dx	=	1	;	Dy	=	-1	;	end
                50	:	begin	Vx	=	9	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	10	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	10	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	6	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
                70	:	begin	Vx	=	6	;	Vy	=	7	;	Dx	=	1	;	Dy	=	-1	;	end
                75	:	begin	Vx	=	9	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	2	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	10	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	5	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
                95	:	begin	Vx	=	7	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                100	:	begin	Vx	=	8	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	3	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	10	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	4	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	-1	;	end
                120	:	begin	Vx	=	8	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                125	:	begin	Vx	=	7	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	4	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	10	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                140	:	begin	Vx	=	2	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	-1	;	end
                145	:	begin	Vx	=	8	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                150	:	begin	Vx	=	6	;	Vy	=	8	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	5	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	10	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                165	:	begin	Vx	=	1	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	-1	;	end
                170	:	begin	Vx	=	9	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                175	:	begin	Vx	=	5	;	Vy	=	9	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	6	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	10	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	9	;	Dx	=	1	;	Dy	=	-1	;	end
                195	:	begin	Vx	=	9	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                200	:	begin	Vx	=	4	;	Vy	=	9	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	7	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	9	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                215	:	begin	Vx	=	1	;	Vy	=	9	;	Dx	=	1	;	Dy	=	-1	;	end
                220	:	begin	Vx	=	9	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                225	:	begin	Vx	=	3	;	Vy	=	10	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	8	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	9	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                240	:	begin	Vx	=	3	;	Vy	=	9	;	Dx	=	1	;	Dy	=	-1	;	end
                245	:	begin	Vx	=	9	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	2	;	Vy	=	10	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	9	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	8	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                265	:	begin	Vx	=	4	;	Vy	=	8	;	Dx	=	1	;	Dy	=	-1	;	end
                270	:	begin	Vx	=	9	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	1	;	Vy	=	10	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	10	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	7	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end
                290	:	begin	Vx	=	5	;	Vy	=	8	;	Dx	=	1	;	Dy	=	-1	;	end
                295	:	begin	Vx	=	9	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	1	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	10	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	6	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
                315	:	begin	Vx	=	6	;	Vy	=	7	;	Dx	=	1	;	Dy	=	-1	;	end
                320	:	begin	Vx	=	9	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	2	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	10	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	5	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	-1	;	end
                340	:	begin	Vx	=	7	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                345	:	begin	Vx	=	8	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	3	;	Vy	=	10	;	Dx	=	-1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	10	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	3	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	-1	;	end

            endcase
            9 : case(deg)
                0	:	begin	Vx	=	9	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	2	;	Vy	=	9	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	8	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	7	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                20	:	begin	Vx	=	3	;	Vy	=	8	;	Dx	=	1	;	Dy	=	-1	;	end
                25	:	begin	Vx	=	8	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	1	;	Vy	=	9	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	9	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	7	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                45	:	begin	Vx	=	4	;	Vy	=	7	;	Dx	=	1	;	Dy	=	-1	;	end
                50	:	begin	Vx	=	8	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	9	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	9	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	6	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end
                70	:	begin	Vx	=	5	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                75	:	begin	Vx	=	8	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	1	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	9	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	5	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
                95	:	begin	Vx	=	6	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                100	:	begin	Vx	=	7	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	3	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	9	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	3	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
                120	:	begin	Vx	=	7	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                125	:	begin	Vx	=	7	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	4	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	9	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                140	:	begin	Vx	=	2	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
                145	:	begin	Vx	=	7	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                150	:	begin	Vx	=	6	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	5	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	9	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                165	:	begin	Vx	=	1	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
                170	:	begin	Vx	=	8	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                175	:	begin	Vx	=	5	;	Vy	=	8	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	6	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	9	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	8	;	Dx	=	1	;	Dy	=	-1	;	end
                195	:	begin	Vx	=	8	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                200	:	begin	Vx	=	4	;	Vy	=	8	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	7	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	8	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                215	:	begin	Vx	=	1	;	Vy	=	8	;	Dx	=	1	;	Dy	=	-1	;	end
                220	:	begin	Vx	=	8	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                225	:	begin	Vx	=	3	;	Vy	=	9	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	8	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	8	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                240	:	begin	Vx	=	2	;	Vy	=	8	;	Dx	=	1	;	Dy	=	-1	;	end
                245	:	begin	Vx	=	8	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	2	;	Vy	=	9	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	8	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	7	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                265	:	begin	Vx	=	4	;	Vy	=	8	;	Dx	=	1	;	Dy	=	-1	;	end
                270	:	begin	Vx	=	8	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	0	;	Vy	=	9	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	9	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	6	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                290	:	begin	Vx	=	5	;	Vy	=	7	;	Dx	=	1	;	Dy	=	-1	;	end
                295	:	begin	Vx	=	8	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	1	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	9	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	5	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end
                315	:	begin	Vx	=	6	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                320	:	begin	Vx	=	8	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	2	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	9	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	4	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
                340	:	begin	Vx	=	6	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                345	:	begin	Vx	=	7	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	3	;	Vy	=	9	;	Dx	=	-1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	9	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	3	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	-1	;	end
            endcase
            8 : case(deg)
                0	:	begin	Vx	=	8	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	2	;	Vy	=	8	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	7	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	7	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                20	:	begin	Vx	=	3	;	Vy	=	7	;	Dx	=	1	;	Dy	=	-1	;	end
                25	:	begin	Vx	=	7	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	1	;	Vy	=	8	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	8	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	6	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                45	:	begin	Vx	=	4	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                50	:	begin	Vx	=	7	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	8	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	8	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	5	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                70	:	begin	Vx	=	5	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                75	:	begin	Vx	=	7	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	1	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	8	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	4	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end
                95	:	begin	Vx	=	5	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                100	:	begin	Vx	=	6	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	2	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	8	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	3	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end
                120	:	begin	Vx	=	6	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                125	:	begin	Vx	=	6	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	3	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	8	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                140	:	begin	Vx	=	2	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end
                145	:	begin	Vx	=	7	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                150	:	begin	Vx	=	5	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	4	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	8	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                165	:	begin	Vx	=	1	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end
                170	:	begin	Vx	=	7	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                175	:	begin	Vx	=	4	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	5	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	8	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	7	;	Dx	=	1	;	Dy	=	-1	;	end
                195	:	begin	Vx	=	7	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                200	:	begin	Vx	=	3	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	6	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	8	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                215	:	begin	Vx	=	1	;	Vy	=	7	;	Dx	=	1	;	Dy	=	-1	;	end
                220	:	begin	Vx	=	7	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                225	:	begin	Vx	=	2	;	Vy	=	8	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	7	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	7	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                240	:	begin	Vx	=	2	;	Vy	=	7	;	Dx	=	1	;	Dy	=	-1	;	end
                245	:	begin	Vx	=	7	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	1	;	Vy	=	8	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	7	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	6	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                265	:	begin	Vx	=	3	;	Vy	=	7	;	Dx	=	1	;	Dy	=	-1	;	end
                270	:	begin	Vx	=	7	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	0	;	Vy	=	8	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	8	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	6	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                290	:	begin	Vx	=	4	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                295	:	begin	Vx	=	7	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	1	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	8	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	5	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                315	:	begin	Vx	=	5	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                320	:	begin	Vx	=	7	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	2	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	8	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	4	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end
                340	:	begin	Vx	=	6	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                345	:	begin	Vx	=	6	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	3	;	Vy	=	8	;	Dx	=	-1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	8	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	3	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	-1	;	end

            endcase
            7 : case(deg)
                0	:	begin	Vx	=	7	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	1	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	6	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	6	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                20	:	begin	Vx	=	2	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                25	:	begin	Vx	=	6	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	1	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	7	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	5	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                45	:	begin	Vx	=	3	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                50	:	begin	Vx	=	6	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	7	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	7	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	4	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                70	:	begin	Vx	=	4	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                75	:	begin	Vx	=	6	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	1	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	7	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	4	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                95	:	begin	Vx	=	5	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                100	:	begin	Vx	=	6	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	2	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	7	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	3	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                120	:	begin	Vx	=	5	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                125	:	begin	Vx	=	5	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	3	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	7	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                140	:	begin	Vx	=	2	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                145	:	begin	Vx	=	6	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                150	:	begin	Vx	=	4	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	4	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	7	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                165	:	begin	Vx	=	1	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                170	:	begin	Vx	=	6	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                175	:	begin	Vx	=	4	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	5	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	7	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                195	:	begin	Vx	=	6	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                200	:	begin	Vx	=	3	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	5	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	7	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                215	:	begin	Vx	=	1	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                220	:	begin	Vx	=	6	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                225	:	begin	Vx	=	2	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	6	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	6	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                240	:	begin	Vx	=	2	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                245	:	begin	Vx	=	6	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	1	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	7	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	6	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                265	:	begin	Vx	=	3	;	Vy	=	6	;	Dx	=	1	;	Dy	=	-1	;	end
                270	:	begin	Vx	=	6	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	0	;	Vy	=	7	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	7	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	5	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                290	:	begin	Vx	=	3	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                295	:	begin	Vx	=	6	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	1	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	7	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	4	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                315	:	begin	Vx	=	4	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                320	:	begin	Vx	=	6	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	2	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	7	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	3	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end
                340	:	begin	Vx	=	5	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                345	:	begin	Vx	=	5	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	2	;	Vy	=	7	;	Dx	=	-1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	7	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	2	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	-1	;	end

            endcase
            6 : case(deg)
                0	:	begin	Vx	=	6	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	1	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	6	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	5	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                20	:	begin	Vx	=	2	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                25	:	begin	Vx	=	5	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	0	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	6	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	5	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                45	:	begin	Vx	=	3	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                50	:	begin	Vx	=	5	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	6	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	6	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	4	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                70	:	begin	Vx	=	3	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                75	:	begin	Vx	=	5	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	1	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	6	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	3	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                95	:	begin	Vx	=	4	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                100	:	begin	Vx	=	5	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	2	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	6	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	2	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                120	:	begin	Vx	=	4	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                125	:	begin	Vx	=	4	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	3	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	6	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                140	:	begin	Vx	=	2	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                145	:	begin	Vx	=	5	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                150	:	begin	Vx	=	4	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	3	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	6	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                165	:	begin	Vx	=	1	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                170	:	begin	Vx	=	5	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                175	:	begin	Vx	=	3	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	4	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	6	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                195	:	begin	Vx	=	5	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                200	:	begin	Vx	=	2	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	5	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	6	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                215	:	begin	Vx	=	1	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                220	:	begin	Vx	=	5	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                225	:	begin	Vx	=	2	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	5	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	5	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                240	:	begin	Vx	=	1	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                245	:	begin	Vx	=	5	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	1	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	6	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	5	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                265	:	begin	Vx	=	2	;	Vy	=	5	;	Dx	=	1	;	Dy	=	-1	;	end
                270	:	begin	Vx	=	5	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	0	;	Vy	=	6	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	6	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	4	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                290	:	begin	Vx	=	3	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                295	:	begin	Vx	=	5	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	1	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	6	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	4	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                315	:	begin	Vx	=	4	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                320	:	begin	Vx	=	5	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	1	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	6	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	3	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end
                340	:	begin	Vx	=	4	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                345	:	begin	Vx	=	5	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	2	;	Vy	=	6	;	Dx	=	-1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	6	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	2	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	-1	;	end

            endcase
            5 : case(deg)
                0	:	begin	Vx	=	5	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	1	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	5	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	4	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                20	:	begin	Vx	=	2	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                25	:	begin	Vx	=	4	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	0	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	5	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	4	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                45	:	begin	Vx	=	2	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                50	:	begin	Vx	=	4	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	5	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	5	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	3	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                70	:	begin	Vx	=	3	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                75	:	begin	Vx	=	4	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	1	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	5	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	3	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                95	:	begin	Vx	=	3	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                100	:	begin	Vx	=	4	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	2	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	5	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	2	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                120	:	begin	Vx	=	4	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                125	:	begin	Vx	=	3	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	2	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	5	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                140	:	begin	Vx	=	1	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                145	:	begin	Vx	=	4	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                150	:	begin	Vx	=	3	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	3	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	5	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                165	:	begin	Vx	=	1	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                170	:	begin	Vx	=	4	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                175	:	begin	Vx	=	2	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	3	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	5	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                195	:	begin	Vx	=	4	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                200	:	begin	Vx	=	2	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	4	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	5	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                215	:	begin	Vx	=	0	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                220	:	begin	Vx	=	4	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                225	:	begin	Vx	=	1	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	4	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	5	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                240	:	begin	Vx	=	1	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                245	:	begin	Vx	=	4	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	1	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	5	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	4	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                265	:	begin	Vx	=	2	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                270	:	begin	Vx	=	4	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	0	;	Vy	=	5	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	5	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	4	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                290	:	begin	Vx	=	2	;	Vy	=	4	;	Dx	=	1	;	Dy	=	-1	;	end
                295	:	begin	Vx	=	4	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	1	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	5	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	3	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                315	:	begin	Vx	=	3	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                320	:	begin	Vx	=	4	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	1	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	5	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	3	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end
                340	:	begin	Vx	=	3	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                345	:	begin	Vx	=	4	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	2	;	Vy	=	5	;	Dx	=	-1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	5	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	2	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	-1	;	end

            endcase
            4 : case(deg)
                0	:	begin	Vx	=	4	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	1	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	4	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	4	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                20	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                25	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	0	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	4	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                45	:	begin	Vx	=	2	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                50	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	4	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	4	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	3	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                70	:	begin	Vx	=	2	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                75	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	1	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	4	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	2	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                95	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                100	:	begin	Vx	=	3	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	1	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	4	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	2	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                120	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                125	:	begin	Vx	=	3	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	2	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	4	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                140	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                145	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                150	:	begin	Vx	=	2	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	2	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	4	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                165	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                170	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                175	:	begin	Vx	=	2	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	3	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	4	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                195	:	begin	Vx	=	3	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                200	:	begin	Vx	=	1	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	3	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	4	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                215	:	begin	Vx	=	0	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                220	:	begin	Vx	=	3	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                225	:	begin	Vx	=	1	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	4	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	4	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                240	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                245	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	0	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	4	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                265	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                270	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	0	;	Vy	=	4	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	4	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	3	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                290	:	begin	Vx	=	2	;	Vy	=	3	;	Dx	=	1	;	Dy	=	-1	;	end
                295	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	1	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	4	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	3	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                315	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                320	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	1	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	4	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	2	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end
                340	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                345	:	begin	Vx	=	3	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	2	;	Vy	=	4	;	Dx	=	-1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	4	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	2	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	-1	;	end

            endcase
            3 : case(deg)
                0	:	begin	Vx	=	3	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	0	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                20	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                25	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	0	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                45	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                50	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	3	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                70	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                75	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                95	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                100	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                120	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                125	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	2	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	3	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                140	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                145	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                150	:	begin	Vx	=	2	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	2	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	3	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                165	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                170	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                175	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	2	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                195	:	begin	Vx	=	2	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                200	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	3	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                215	:	begin	Vx	=	0	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                220	:	begin	Vx	=	2	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                225	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                240	:	begin	Vx	=	0	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                245	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	0	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                265	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                270	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	0	;	Vy	=	3	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	3	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                290	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                295	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                315	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	1	;	Dy	=	-1	;	end
                320	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
                340	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                345	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	1	;	Vy	=	3	;	Dx	=	-1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	3	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	-1	;	end
            endcase
            2 : case(deg)
                0	:	begin	Vx	=	2	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	0	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                20	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                25	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	0	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                45	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                50	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	2	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                70	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                75	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                95	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                100	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                120	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                125	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	2	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                140	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                145	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                150	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	2	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                165	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                170	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                175	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	2	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                195	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                200	:	begin	Vx	=	0	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	2	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                215	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                220	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                225	:	begin	Vx	=	0	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                240	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                245	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	0	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	2	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                265	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                270	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	0	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                290	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                295	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                315	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                320	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
                340	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	1	;	Dy	=	-1	;	end
                345	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	1	;	Vy	=	2	;	Dx	=	-1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	2	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	-1	;	end
            endcase
            1 : case(deg)
                0	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                20	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                25	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                45	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                50	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                70	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                75	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                95	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                100	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                120	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                125	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                140	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                145	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                150	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                165	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                170	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                175	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                195	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                200	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                215	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                220	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                225	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                240	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                245	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                265	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                270	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                290	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                295	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                315	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                320	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
                340	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                345	:	begin	Vx	=	0	;	Vy	=	1	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	1	;	Vy	=	1	;	Dx	=	-1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	1	;	Vy	=	0	;	Dx	=	-1	;	Dy	=	1	;	end
            endcase
            0 : case(deg)
                0	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                5	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                10	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                15	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                20	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                25	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                30	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                35	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                40	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                45	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                50	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                55	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	0	;	Dy	=	1	;	end
                60	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                65	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                70	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                75	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                80	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                85	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                90	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                95	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                100	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                105	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                110	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                115	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                120	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                125	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                130	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                135	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                140	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                145	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                150	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                155	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                160	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                165	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                170	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                175	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                180	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                185	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                190	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                195	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                200	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                205	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                210	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                215	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                220	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                225	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                230	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                235	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                240	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                245	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                250	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                255	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                260	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                265	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                270	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                275	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                280	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                285	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                290	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                295	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                300	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                305	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                310	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                315	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                320	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                325	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                330	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                335	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                340	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                345	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                350	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                355	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
                360	:	begin	Vx	=	0	;	Vy	=	0	;	Dx	=	1	;	Dy	=	1	;	end
            endcase
        endcase
    end
end